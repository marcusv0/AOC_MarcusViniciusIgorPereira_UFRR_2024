LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DIV_INSTRUCAO IS
    PORT(
        INSTRUCTION     : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        OPCODE, ADDRESS : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        RS,RT           : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
    );
END DIV_INSTRUCAO;

ARCHITECTURE BEHAVIOR OF DIV_INSTRUCAO IS
BEGIN
    OPCODE <= INSTRUCTION(7 DOWNTO 4);
    RS <= INSTRUCTION(3 DOWNTO 2);
    RT <= INSTRUCTION(1 DOWNTO 0);
    ADDRESS <= INSTRUCTION(3 DOWNTO 0);
END;